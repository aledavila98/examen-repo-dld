`define ADD 4'd0
`define SUB 4'd1
`define MUL 4'd2
`define DIV 4'd3
`define MOD 4'd4
`define AND 4'd5
`define OR  4'd6
`define XOR 4'd7
`define NOT 4'd8
`define SHL 4'd9
`define SHR 4'd10
`define SLT 4'd11
`define SLTU 4'd12
